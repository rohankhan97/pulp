module tb;

endmodule
