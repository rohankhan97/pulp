class cpi_sequencer extends uvm_sequencer#(cpi_frame_item);
	`uvm_component_utils(cpi_sequencer)
	`uvm_component_new
endclass : cpi_sequencer