`define TLM_MASTER