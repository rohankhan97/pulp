//-----------------------------------------------------------------------------
// Title         : Sequence Item Type for Virtual Stdout Monitor
//-----------------------------------------------------------------------------
// File          : vstdout_seq_item.sv
// Author        : Manuel Eggimann  <meggimann@iis.ee.ethz.ch>
// Created       : 08.10.2021
//-----------------------------------------------------------------------------
// Description :
//
// This class implements the primitive sequence item generated by the virtual
// stdout monitor.
//
//-----------------------------------------------------------------------------
// Copyright (C) 2021 ETH Zurich, University of Bologna
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License. You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.
// SPDX-License-Identifier: SHL-0.51
//-----------------------------------------------------------------------------

class vstdout_seq_item extends uvm_sequence_item;
  string channel_name;
  string message;

  `uvm_object_utils_begin(vstdout_seq_item)
    `uvm_field_string(channel_name, UVM_DEFAULT)
    `uvm_field_string(message, UVM_DEFAULT)
  `uvm_object_utils_end
  `uvm_object_new
endclass
