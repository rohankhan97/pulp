package qvip_env_pkg;
	import mgc_i3c_pkg::*;
  import mgc_spi_v1_0_pkg::*;
endpackage
